module hulf_adder (a, b, cout, sum);
    input a, b;
    output cout, sum;

    assign sum = a ^ b;  // XOR for sum
    assign cout = a & b; // AND for carry out

endmodule
